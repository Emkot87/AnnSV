import ann_pkg::*;

module layer(

);



endmodule