package ann_pkg;
    parameter int neuron_size = 8;
    parameter int word_size   = 32;
endpackage