
module ann(
    input 
);

    //layer 1

    genvar i;
    generate
        for 
    endgenerate

    neuron i_neuron(
        
    );

    ram i_ram(

    );

    apb_slave i_apb(

    );

endmodule