module ram(

);

endmodule